module ObjColision(

    );

endmodule