module ObjColision(
        
    );

endmodule